module Register_File (
    input clk, WE3, rst,
    input [4:0] A1, A2, A3,
    input [31:0] WD3,
    output [31:0] RD1, RD2
);
    reg [31:0] reg_mem [31:0];

    integer i;
    always @(posedge clk or negedge rst) begin
        if (!rst) begin
            for(i=0; i<32; i=i+1) begin 
                reg_mem[i] <= 32'd0;
            end

        end
        
        else if(WE3) begin
            reg_mem[A3] <= WD3;
        end
    end

    assign RD1 = (A1 != 0) ? reg_mem[A1] : 0;
    assign RD2 = (A2 != 0) ? reg_mem[A2] : 0;

endmodule